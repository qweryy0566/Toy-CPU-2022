`include "config.v"

module ICache (

);

endmodule